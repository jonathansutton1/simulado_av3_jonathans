-- Elementos de Sistemas
-- developed by Luciano Soares
-- file: Q2_ControlUnit.vhd
-- date: 4/4/2017
-- Modificação:
--   - Rafael Corsi : nova versão: adicionado reg S
--
-- Unidade que controla os componentes da CPU

library ieee;
use ieee.std_logic_1164.all;

entity Q2_ControlUnit is
    port(
		instruction                 : in STD_LOGIC_VECTOR(17 downto 0);  -- instrução para executar
		zr,ng                       : in STD_LOGIC;                      -- valores zr(se zero) e
                                                                     -- ng (se negativo) da ALU
		muxALUI_A                   : out STD_LOGIC;                     -- mux que seleciona entre
                                                                     -- instrução  e ALU para reg. A
		muxAM                       : out STD_LOGIC;                     -- mux que seleciona entre
		zx, nx, zy, ny, f, no       : out STD_LOGIC;                     -- sinais de controle da ALU
		loadA, loadD, loadM, loadPC : out STD_LOGIC               -- sinais de load do reg. A,
                                                                     -- reg. D, Mem. RAM e Program Counter
    );
end entity;

architecture arch of Q2_ControlUnit is

signal jg : std_logic;

begin

  loadPC <= jg and instruction(17) and instruction(0);

  -- implementar somente o loadD para o caso do jgu e jgs
  jg <= '1' when instruction(16) = '0' and ng = '0' and zr = '0' else
        '1' when instruction(16) = '1' and zr = '0' else
        '0';

end architecture;
